// Copyright goes here ;)
// Top.v just top level for proper pinout.

module top (
input wire clk;
input wire reset;
output wire [3:0] dac_out;
)


endmodule
